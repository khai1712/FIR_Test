module Filter_block_1
#(
    parameter n = 63,
    parameter signed [0:16*n-1] coef = 
    {
    16'b1111111111111111,
    16'b1111111111111111,
    16'b1111111111111111,
    16'b1111111111111110,
    16'b1111111111111110,
    16'b1111111111111110,
    16'b1111111111111111,
    16'b0000000000000000,
    16'b0000000000000001,
    16'b0000000000000010,
    16'b0000000000000100,
    16'b0000000000000101,
    16'b0000000000000101,
    16'b0000000000000101,
    16'b0000000000000011,
    16'b1111111111111111,
    16'b1111111111111011,
    16'b1111111111110110,
    16'b1111111111110001,
    16'b1111111111101101,
    16'b1111111111101100,
    16'b1111111111101110,
    16'b1111111111110100,
    16'b0000000000000000,
    16'b0000000000001111,
    16'b0000000000100010,
    16'b0000000000110111,
    16'b0000000001001100,
    16'b0000000001100000,
    16'b0000000001101111,
    16'b0000000001111001,
    16'b0000000001111101,
    16'b0000000001111001,
    16'b0000000001101111,
    16'b0000000001100000,
    16'b0000000001001100,
    16'b0000000000110111,
    16'b0000000000100010,
    16'b0000000000001111,
    16'b0000000000000000,
    16'b1111111111110100,
    16'b1111111111101110,
    16'b1111111111101100,
    16'b1111111111101101,
    16'b1111111111110001,
    16'b1111111111110110,
    16'b1111111111111011,
    16'b1111111111111111,
    16'b0000000000000011,
    16'b0000000000000101,
    16'b0000000000000101,
    16'b0000000000000101,
    16'b0000000000000100,
    16'b0000000000000010,
    16'b0000000000000001,
    16'b0000000000000000,
    16'b1111111111111111,
    16'b1111111111111110,
    16'b1111111111111110,
    16'b1111111111111110,
    16'b1111111111111111,
    16'b1111111111111111,
    16'b1111111111111111
    }
)

(
    input clk, 
    input rst_p, 
    input signed [15:0] x_in,
    input signed [15:0] y_in,
    output reg signed [15:0] x_out,
    output reg signed [15:0] y_out
);  
    reg [15:0] mul;
    reg signed [0:16*(n-1)-1] delay_x;
    integer i, j, k;
    reg signed [15:0] sum;
    
    //for(l=0; l<n; l=l+1) begin
    //    coef_cov[16*k +: 16] = (coef[16*l] == 1'b1) ? {8'b11111111, coef[16*l +: 16]} : {8'b00000000, coef[16*l +: 16]};
    //end

    always @(posedge clk or posedge rst_p) begin
        if(rst_p) begin
            for(i=0; i<n-1; i=i+1) begin
                delay_x[16*i +: 16] <= 0;
            end
            //sum <= 0; 
            x_out <= 0;
            //y_out <= 0;
        end
        else begin
            delay_x[0:15] <= x_in;
            x_out <= delay_x[16*(n-2):16*(n-1)-1];
            for(j=1; j<n-1; j=j+1) begin
                delay_x[16*j +: 16] <= delay_x[16*(j-1) +: 16];
            end
        end
    end
    
    always @(x_in or delay_x) begin
        sum = 0;
        mul = (x_in) * (coef[0:15]); //Lấy 16 bit cuối của phép nhân
        sum = sum + mul; 
        for(k=0; k<n-1; k=k+1) begin
            mul = delay_x[16*k +: 16] * coef[16*(k+1) +: 16];
            sum = sum + mul; //Lấy 16 bit cuối của phép nhân
        end
    end
    
    always @(posedge clk) begin
        y_out <= sum;
    end

endmodule